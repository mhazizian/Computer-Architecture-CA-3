// ALU Functions

`define ADD_FN 3'b000
`define ADDC_FN 3'b001
`define SUB_FN 3'b010
`define SUBC_FN 3'b011
`define AND_FN 3'b100
`define OR_FN 3'b101
